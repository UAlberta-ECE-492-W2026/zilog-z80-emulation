
`timescale 1ns/1ps
`include "alu_op.sv"

module datapath (
    input logic clk,
    input logic reset,

    


)
endmodule
// ###########################
// End of module datapath
// ###########################
